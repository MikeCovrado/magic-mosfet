magic
tech sky130A
timestamp 1610746791
<< nmos >>
rect 35 -5 50 60
<< ndiff >>
rect -25 40 35 60
rect -25 15 -10 40
rect 15 15 35 40
rect -25 -5 35 15
rect 50 40 110 60
rect 50 15 70 40
rect 95 15 110 40
rect 50 -5 110 15
<< ndiffc >>
rect -10 15 15 40
rect 70 15 95 40
<< poly >>
rect 35 60 50 100
rect 35 -25 50 -5
rect -5 -35 50 -25
rect -5 -60 10 -35
rect 35 -60 50 -35
rect -5 -70 50 -60
<< polycont >>
rect 10 -60 35 -35
<< locali >>
rect -50 40 25 50
rect -50 37 -10 40
rect -50 20 -45 37
rect -28 20 -10 37
rect -50 15 -10 20
rect 15 15 25 40
rect -50 5 25 15
rect 60 45 135 50
rect 60 40 170 45
rect 60 15 70 40
rect 95 20 114 40
rect 132 20 170 40
rect 95 15 170 20
rect 60 12 170 15
rect 60 5 135 12
rect -35 -35 45 -25
rect -15 -60 10 -35
rect 35 -60 45 -35
rect -35 -70 45 -60
<< viali >>
rect -45 20 -28 37
rect 114 20 132 40
rect -35 -60 -15 -35
<< metal1 >>
rect -87 37 -20 45
rect -87 20 -45 37
rect -28 20 -20 37
rect -87 13 -20 20
rect 105 40 170 45
rect 105 20 114 40
rect 132 20 170 40
rect 105 12 170 20
rect -80 -35 -5 -25
rect -80 -60 -35 -35
rect -15 -60 -5 -35
rect -80 -70 -5 -60
<< labels >>
rlabel metal1 -80 20 -60 40 1 source
rlabel metal1 145 20 165 40 1 drain
rlabel metal1 -70 -56 -50 -36 1 gate
<< end >>
